library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GFX1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GFX1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"9C",X"63",X"41",X"9C",X"BE",X"BE",X"41",X"00",X"41",X"14",X"36",X"41",X"63",X"63",X"14",X"00",
		X"41",X"41",X"FF",X"00",X"41",X"41",X"FF",X"00",X"00",X"22",X"77",X"00",X"00",X"00",X"77",X"00",
		X"41",X"FF",X"DD",X"63",X"C9",X"77",X"DD",X"00",X"63",X"14",X"55",X"22",X"77",X"36",X"14",X"00",
		X"36",X"C9",X"C9",X"22",X"FF",X"63",X"C9",X"00",X"14",X"14",X"77",X"00",X"36",X"14",X"55",X"00",
		X"14",X"14",X"FF",X"9C",X"FF",X"9C",X"14",X"00",X"00",X"63",X"77",X"00",X"77",X"41",X"36",X"00",
		X"BE",X"41",X"41",X"22",X"FF",X"63",X"41",X"00",X"00",X"55",X"55",X"77",X"55",X"77",X"55",X"00",
		X"36",X"C9",X"C9",X"BE",X"FF",X"FF",X"C9",X"00",X"00",X"36",X"14",X"41",X"14",X"63",X"14",X"00",
		X"00",X"77",X"88",X"00",X"00",X"00",X"FF",X"00",X"36",X"14",X"55",X"36",X"77",X"36",X"14",X"00",
		X"36",X"C9",X"DD",X"36",X"77",X"C9",X"DD",X"00",X"00",X"55",X"14",X"63",X"63",X"77",X"14",X"00",
		X"9C",X"C9",X"EB",X"00",X"BE",X"C9",X"C9",X"00",X"63",X"14",X"14",X"63",X"77",X"77",X"14",X"00",
		X"62",X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"41",X"00",X"00",X"00",X"62",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"94",
		X"62",X"62",X"63",X"63",X"63",X"63",X"62",X"62",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"94",X"94",X"9C",X"9C",X"9C",X"9C",X"94",X"94",
		X"F6",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F6",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F6",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F6",
		X"08",X"01",X"02",X"0C",X"0C",X"02",X"01",X"08",X"01",X"08",X"04",X"03",X"03",X"04",X"08",X"01",
		X"08",X"81",X"02",X"0C",X"0C",X"02",X"81",X"08",X"01",X"48",X"04",X"03",X"03",X"04",X"48",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"08",X"31",X"9A",X"84",X"84",X"9A",X"31",X"08",X"01",X"38",X"65",X"42",X"42",X"65",X"38",X"01",
		X"9C",X"4F",X"B1",X"2E",X"B2",X"4F",X"4F",X"9C",X"63",X"8F",X"F8",X"17",X"74",X"8F",X"8F",X"63",
		X"9C",X"F1",X"4F",X"2E",X"2E",X"4F",X"F1",X"9C",X"63",X"F8",X"8F",X"17",X"17",X"8F",X"F8",X"63",
		X"9C",X"4F",X"4F",X"B2",X"2E",X"F1",X"4F",X"9C",X"63",X"8F",X"8F",X"74",X"17",X"F8",X"8F",X"63",
		X"00",X"84",X"08",X"00",X"00",X"08",X"84",X"00",X"00",X"42",X"01",X"00",X"00",X"01",X"42",X"00",
		X"00",X"86",X"08",X"08",X"08",X"08",X"86",X"00",X"00",X"46",X"01",X"01",X"01",X"01",X"46",X"00",
		X"08",X"87",X"08",X"08",X"08",X"08",X"87",X"08",X"01",X"4E",X"01",X"01",X"01",X"01",X"4E",X"01",
		X"02",X"C8",X"04",X"22",X"02",X"14",X"78",X"22",X"14",X"B1",X"22",X"04",X"14",X"02",X"C1",X"04",
		X"20",X"49",X"10",X"02",X"20",X"04",X"F7",X"02",X"04",X"FE",X"02",X"10",X"04",X"20",X"89",X"10",
		X"22",X"81",X"14",X"20",X"22",X"10",X"8F",X"20",X"10",X"4F",X"20",X"14",X"10",X"22",X"48",X"14",
		X"08",X"B1",X"92",X"84",X"84",X"92",X"B1",X"08",X"01",X"78",X"64",X"42",X"42",X"64",X"78",X"01",
		X"00",X"92",X"84",X"08",X"08",X"84",X"92",X"00",X"00",X"64",X"42",X"01",X"01",X"42",X"64",X"00",
		X"00",X"84",X"08",X"00",X"00",X"08",X"84",X"00",X"00",X"42",X"01",X"00",X"00",X"01",X"42",X"00",
		X"00",X"04",X"08",X"00",X"00",X"08",X"04",X"00",X"00",X"02",X"01",X"00",X"00",X"01",X"02",X"00",
		X"00",X"02",X"04",X"08",X"08",X"04",X"02",X"00",X"00",X"04",X"02",X"01",X"01",X"02",X"04",X"00",
		X"08",X"01",X"02",X"04",X"04",X"02",X"01",X"08",X"01",X"08",X"04",X"02",X"02",X"04",X"08",X"01",
		X"08",X"B1",X"92",X"84",X"84",X"92",X"B1",X"08",X"01",X"78",X"64",X"42",X"42",X"64",X"78",X"01",
		X"08",X"B1",X"9E",X"8C",X"8C",X"9E",X"B1",X"08",X"01",X"78",X"67",X"43",X"43",X"67",X"78",X"01",
		X"08",X"BF",X"92",X"84",X"84",X"92",X"BF",X"08",X"01",X"7F",X"64",X"42",X"42",X"64",X"7F",X"01",
		X"0C",X"B9",X"B1",X"92",X"92",X"B1",X"B9",X"0C",X"03",X"79",X"78",X"64",X"64",X"78",X"79",X"03",
		X"0C",X"B5",X"BD",X"92",X"92",X"BD",X"B5",X"0C",X"03",X"7A",X"7B",X"64",X"64",X"7B",X"7A",X"03",
		X"0C",X"B3",X"B3",X"9E",X"9E",X"B3",X"B3",X"0C",X"03",X"7C",X"7C",X"67",X"67",X"7C",X"7C",X"03",
		X"00",X"00",X"36",X"36",X"36",X"36",X"00",X"00",X"00",X"00",X"36",X"36",X"36",X"36",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"88",X"36",X"22",X"88",X"9C",X"9C",X"22",X"00",X"63",X"88",X"9C",X"63",X"77",X"77",X"88",X"00",
		X"22",X"22",X"BE",X"00",X"22",X"22",X"BE",X"00",X"00",X"14",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"22",X"BE",X"AA",X"36",X"22",X"BE",X"AA",X"00",X"36",X"C9",X"EB",X"14",X"FF",X"9C",X"C9",X"00",
		X"9C",X"22",X"22",X"14",X"BE",X"36",X"22",X"00",X"88",X"C9",X"FF",X"00",X"DD",X"88",X"EB",X"00",
		X"88",X"88",X"BE",X"88",X"BE",X"88",X"88",X"00",X"00",X"36",X"FF",X"41",X"FF",X"63",X"9C",X"00",
		X"9C",X"22",X"22",X"14",X"BE",X"36",X"22",X"00",X"41",X"AA",X"AA",X"BE",X"EB",X"BE",X"AA",X"00",
		X"9C",X"22",X"22",X"9C",X"BE",X"BE",X"22",X"00",X"00",X"DD",X"C9",X"63",X"C9",X"77",X"C9",X"00",
		X"00",X"BE",X"00",X"00",X"00",X"00",X"BE",X"00",X"9C",X"88",X"EB",X"9C",X"BE",X"9C",X"C9",X"00",
		X"9C",X"22",X"AA",X"9C",X"BE",X"22",X"AA",X"00",X"00",X"EB",X"C9",X"36",X"36",X"FF",X"C9",X"00",
		X"88",X"22",X"36",X"00",X"9C",X"22",X"22",X"00",X"77",X"C9",X"C9",X"36",X"FF",X"FF",X"C9",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BE",X"88",X"88",X"BE",X"BE",X"BE",X"88",X"00",X"63",X"9C",X"9C",X"63",X"77",X"77",X"88",X"00",
		X"9C",X"22",X"22",X"BE",X"BE",X"BE",X"22",X"00",X"36",X"C9",X"C9",X"FF",X"FF",X"FF",X"C9",X"00",
		X"14",X"36",X"22",X"88",X"36",X"9C",X"22",X"00",X"14",X"9C",X"88",X"63",X"9C",X"77",X"88",X"00",
		X"88",X"22",X"36",X"BE",X"9C",X"BE",X"22",X"00",X"63",X"88",X"9C",X"FF",X"77",X"FF",X"88",X"00",
		X"22",X"BE",X"22",X"00",X"22",X"BE",X"22",X"00",X"88",X"FF",X"C9",X"00",X"C9",X"FF",X"C9",X"00",
		X"00",X"00",X"00",X"BE",X"00",X"BE",X"00",X"00",X"88",X"C9",X"C9",X"FF",X"C9",X"FF",X"C9",X"00",
		X"BE",X"36",X"22",X"88",X"BE",X"9C",X"22",X"00",X"C9",X"9C",X"C9",X"63",X"C9",X"77",X"88",X"00",
		X"BE",X"00",X"00",X"BE",X"BE",X"BE",X"00",X"00",X"FF",X"41",X"41",X"FF",X"FF",X"FF",X"41",X"00",
		X"22",X"22",X"BE",X"00",X"22",X"22",X"BE",X"00",X"88",X"88",X"FF",X"00",X"88",X"88",X"FF",X"00",
		X"9C",X"22",X"22",X"14",X"BE",X"36",X"22",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"22",X"88",X"BE",X"BE",X"36",X"BE",X"9C",X"00",X"88",X"41",X"36",X"FF",X"9C",X"FF",X"63",X"00",
		X"22",X"BE",X"22",X"00",X"22",X"BE",X"22",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"BE",X"00",X"00",X"BE",X"BE",X"BE",X"88",X"00",X"FF",X"77",X"77",X"FF",X"FF",X"FF",X"63",X"00",
		X"BE",X"00",X"9C",X"BE",X"BE",X"BE",X"88",X"00",X"FF",X"77",X"41",X"FF",X"FF",X"FF",X"63",X"00",
		X"9C",X"22",X"22",X"9C",X"BE",X"BE",X"22",X"00",X"77",X"88",X"88",X"77",X"FF",X"FF",X"88",X"00",
		X"00",X"88",X"88",X"BE",X"88",X"BE",X"88",X"00",X"77",X"88",X"88",X"FF",X"FF",X"FF",X"88",X"00",
		X"AA",X"22",X"BE",X"9C",X"9C",X"BE",X"AA",X"00",X"77",X"88",X"88",X"77",X"FF",X"FF",X"88",X"00",
		X"22",X"88",X"BE",X"BE",X"36",X"BE",X"9C",X"00",X"77",X"88",X"C9",X"FF",X"FF",X"FF",X"88",X"00",
		X"9C",X"22",X"22",X"14",X"BE",X"36",X"22",X"00",X"00",X"C9",X"DD",X"36",X"55",X"FF",X"C9",X"00",
		X"00",X"00",X"BE",X"00",X"00",X"00",X"BE",X"00",X"88",X"88",X"FF",X"00",X"88",X"88",X"FF",X"00",
		X"9C",X"22",X"22",X"9C",X"BE",X"BE",X"22",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"9C",X"9C",X"00",X"88",X"88",X"BE",X"00",X"FF",X"41",X"41",X"FF",X"FF",X"FF",X"00",X"00",
		X"BE",X"9C",X"9C",X"BE",X"BE",X"BE",X"88",X"00",X"FF",X"41",X"41",X"FF",X"FF",X"FF",X"63",X"00",
		X"36",X"9C",X"9C",X"36",X"BE",X"BE",X"88",X"00",X"9C",X"77",X"77",X"9C",X"BE",X"BE",X"63",X"00",
		X"00",X"00",X"BE",X"00",X"00",X"00",X"BE",X"00",X"BE",X"FF",X"41",X"00",X"FF",X"BE",X"41",X"00",
		X"22",X"BE",X"22",X"36",X"22",X"BE",X"AA",X"00",X"9C",X"C9",X"FF",X"88",X"BE",X"88",X"EB",X"00",
		X"BD",X"50",X"4A",X"18",X"C8",X"09",X"90",X"50",X"41",X"27",X"50",X"4E",X"19",X"00",X"01",X"00",
		X"BD",X"50",X"4A",X"D8",X"C8",X"09",X"90",X"37",X"41",X"27",X"37",X"4E",X"D9",X"00",X"01",X"00",
		X"BD",X"50",X"4A",X"10",X"C8",X"09",X"90",X"50",X"41",X"67",X"50",X"4E",X"11",X"00",X"01",X"00",
		X"BD",X"34",X"09",X"53",X"C8",X"41",X"52",X"34",X"01",X"FF",X"00",X"C8",X"37",X"BD",X"4E",X"09",
		X"00",X"88",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"41",X"00",X"00",X"00",X"00",X"41",X"00",
		X"9C",X"22",X"01",X"22",X"22",X"41",X"1C",X"9C",X"63",X"23",X"88",X"14",X"14",X"08",X"14",X"63",
		X"4C",X"47",X"B5",X"4A",X"0B",X"7E",X"C5",X"B8",X"34",X"09",X"9E",X"0A",X"78",X"DC",X"48",X"B5",
		X"C5",X"34",X"0A",X"9E",X"47",X"78",X"B9",X"48",X"B3",X"B3",X"B3",X"B3",X"6F",X"6F",X"6F",X"6F",
		X"9E",X"02",X"63",X"00",X"00",X"90",X"04",X"67",X"00",X"22",X"22",X"00",X"41",X"63",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"9C",X"88",X"00",X"14",X"14",X"00",
		X"10",X"92",X"C8",X"41",X"BD",X"17",X"09",X"93",X"17",X"4E",X"64",X"BD",X"01",X"01",X"00",X"C8",
		X"4A",X"9A",X"50",X"41",X"90",X"17",X"09",X"9B",X"17",X"4E",X"64",X"BD",X"01",X"05",X"00",X"C8",
		X"02",X"88",X"C9",X"55",X"14",X"88",X"89",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"89",X"41",X"22",X"AA",X"C9",X"41",X"04",
		X"00",X"FC",X"C8",X"41",X"BD",X"34",X"09",X"DA",X"13",X"09",X"05",X"10",X"B5",X"02",X"42",X"41",
		X"03",X"00",X"01",X"10",X"10",X"4E",X"6C",X"BD",X"C8",X"09",X"90",X"14",X"4A",X"02",X"50",X"41",
		X"00",X"22",X"00",X"41",X"00",X"22",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"14",X"00",X"88",X"00",X"14",X"00",X"FF",X"86",X"88",X"41",X"88",X"41",X"8A",X"FF",
		X"06",X"AF",X"BD",X"24",X"00",X"4A",X"C8",X"10",X"6A",X"00",X"34",X"23",X"99",X"08",X"FE",X"09",
		X"F1",X"10",X"41",X"21",X"67",X"01",X"24",X"00",X"BD",X"50",X"4A",X"12",X"C8",X"09",X"90",X"35",
		X"41",X"FF",X"35",X"4E",X"13",X"00",X"01",X"00",X"BD",X"62",X"09",X"73",X"C8",X"0A",X"5B",X"35",
		X"0A",X"72",X"35",X"0A",X"13",X"35",X"09",X"32",X"35",X"0A",X"8D",X"35",X"09",X"5E",X"62",X"0A",
		X"76",X"35",X"09",X"1D",X"35",X"0A",X"5D",X"35",X"09",X"C1",X"62",X"0A",X"D7",X"35",X"0A",X"79",
		X"35",X"0A",X"C0",X"35",X"09",X"80",X"35",X"09",X"21",X"35",X"0A",X"C4",X"63",X"0A",X"AC",X"35",
		X"00",X"FF",X"1C",X"89",X"00",X"41",X"00",X"41",X"00",X"88",X"63",X"88",X"00",X"89",X"14",X"FF",
		X"22",X"00",X"00",X"00",X"9C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"35",X"09",X"D1",X"63",X"0A",X"E7",X"35",X"0A",X"FD",X"35",X"0A",X"FC",X"35",X"09",X"9D",X"35",
		X"0A",X"D1",X"35",X"0A",X"BC",X"63",X"09",X"60",X"36",X"09",X"00",X"36",X"0A",X"47",X"36",X"0A",
		X"00",X"14",X"00",X"41",X"00",X"AA",X"00",X"41",X"00",X"02",X"00",X"C9",X"00",X"14",X"00",X"89",
		X"49",X"00",X"22",X"00",X"C9",X"00",X"04",X"00",X"88",X"00",X"55",X"00",X"88",X"00",X"22",X"00",
		X"34",X"BE",X"00",X"09",X"FE",X"23",X"92",X"F3",X"34",X"4A",X"8E",X"50",X"B3",X"01",X"AF",X"09",
		X"F4",X"B5",X"B3",X"47",X"34",X"BF",X"86",X"4A",X"90",X"B5",X"6E",X"46",X"50",X"9A",X"10",X"6E",
		X"00",X"00",X"00",X"9C",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"63",X"00",X"00",X"00",X"22",
		X"41",X"14",X"15",X"00",X"49",X"9C",X"14",X"00",X"22",X"14",X"81",X"00",X"2A",X"63",X"88",X"00",
		X"B5",X"65",X"47",X"09",X"D0",X"17",X"41",X"B6",X"20",X"04",X"01",X"D0",X"6E",X"B5",X"06",X"47",
		X"41",X"B7",X"14",X"6E",X"A2",X"20",X"09",X"01",X"06",X"47",X"B5",X"0E",X"04",X"41",X"D0",X"16",
		X"09",X"01",X"20",X"04",X"D4",X"06",X"6E",X"B5",X"D0",X"14",X"41",X"D6",X"47",X"09",X"9F",X"20",
		X"6E",X"B5",X"06",X"47",X"01",X"D0",X"04",X"41",X"A9",X"20",X"09",X"01",X"16",X"6E",X"D1",X"06",
		X"04",X"41",X"D0",X"15",X"B5",X"A3",X"47",X"09",X"D0",X"06",X"6E",X"B5",X"20",X"04",X"01",X"D0",
		X"47",X"09",X"34",X"20",X"41",X"D5",X"17",X"6E",X"01",X"D0",X"04",X"41",X"06",X"47",X"B5",X"25",
		X"16",X"6E",X"B6",X"06",X"09",X"01",X"20",X"04",X"B5",X"3E",X"47",X"09",X"D0",X"14",X"41",X"D6",
		X"20",X"04",X"01",X"D0",X"6E",X"B5",X"06",X"47",X"41",X"D3",X"16",X"6E",X"B7",X"20",X"09",X"01",
		X"06",X"47",X"B5",X"37",X"04",X"41",X"D0",X"15",X"09",X"01",X"20",X"04",X"D2",X"06",X"6E",X"B5",
		X"D0",X"16",X"41",X"B5",X"47",X"09",X"49",X"20",X"6E",X"B5",X"06",X"47",X"01",X"D0",X"04",X"41",
		X"52",X"20",X"09",X"01",X"15",X"6E",X"B6",X"06",X"04",X"41",X"D0",X"17",X"B5",X"43",X"47",X"09",
		X"D4",X"06",X"6E",X"B5",X"20",X"04",X"01",X"D0",X"47",X"09",X"D4",X"20",X"41",X"D2",X"14",X"6E",
		X"01",X"D0",X"04",X"41",X"06",X"47",X"B5",X"45",X"16",X"6E",X"B5",X"06",X"09",X"01",X"20",X"04",
		X"B5",X"E8",X"47",X"09",X"D0",X"16",X"41",X"D3",X"20",X"04",X"01",X"D0",X"6E",X"B5",X"06",X"47",
		X"41",X"D5",X"15",X"6E",X"E0",X"20",X"09",X"01",X"06",X"47",X"B5",X"72",X"04",X"41",X"D0",X"17",
		X"09",X"01",X"20",X"04",X"B7",X"06",X"6E",X"B5",X"D0",X"20",X"93",X"03",X"47",X"01",X"F3",X"05",
		X"07",X"40",X"26",X"66",X"21",X"60",X"27",X"42",X"03",X"37",X"07",X"09",X"05",X"11",X"41",X"93",
		X"08",X"04",X"01",X"EA",X"6E",X"B5",X"06",X"47",X"6E",X"47",X"B5",X"0E",X"20",X"41",X"80",X"12",
		X"09",X"01",X"08",X"04",X"93",X"06",X"6E",X"B5",X"EA",X"B5",X"6E",X"47",X"47",X"80",X"20",X"41",
		X"B7",X"08",X"09",X"01",X"12",X"6E",X"93",X"06",X"04",X"6E",X"EA",X"B5",X"B5",X"20",X"47",X"80",
		X"47",X"09",X"A2",X"08",X"41",X"93",X"10",X"6E",X"01",X"EA",X"04",X"6E",X"06",X"47",X"B5",X"20",
		X"B5",X"45",X"47",X"09",X"80",X"12",X"41",X"93",X"08",X"04",X"01",X"EA",X"6E",X"B5",X"06",X"47",
		X"6E",X"47",X"B5",X"65",X"20",X"41",X"80",X"13",X"09",X"01",X"08",X"04",X"93",X"06",X"6E",X"B5",
		X"EA",X"B5",X"6E",X"47",X"47",X"80",X"20",X"41",X"D4",X"08",X"09",X"01",X"10",X"6E",X"93",X"06",
		X"04",X"6E",X"EA",X"B5",X"B5",X"20",X"47",X"80",X"47",X"09",X"A9",X"08",X"41",X"93",X"12",X"6E",
		X"01",X"EA",X"04",X"6E",X"06",X"47",X"B5",X"20",X"B5",X"72",X"47",X"09",X"80",X"13",X"41",X"93",
		X"08",X"04",X"01",X"EA",X"6E",X"B5",X"06",X"47",X"6E",X"47",X"B5",X"5F",X"20",X"41",X"80",X"10",
		X"09",X"01",X"08",X"04",X"93",X"06",X"6E",X"B5",X"EA",X"B5",X"6E",X"47",X"47",X"80",X"20",X"41",
		X"A3",X"08",X"09",X"01",X"11",X"6E",X"93",X"06",X"04",X"6E",X"EA",X"B5",X"B5",X"20",X"47",X"80",
		X"47",X"09",X"34",X"08",X"41",X"93",X"13",X"6E",X"01",X"EA",X"04",X"6E",X"06",X"47",X"B5",X"20",
		X"B5",X"25",X"47",X"09",X"80",X"12",X"41",X"93",X"08",X"04",X"01",X"EA",X"6E",X"B5",X"06",X"47",
		X"6E",X"47",X"B5",X"E8",X"20",X"41",X"80",X"12",X"09",X"01",X"08",X"04",X"93",X"06",X"6E",X"B5",
		X"EA",X"B5",X"6E",X"47",X"47",X"80",X"20",X"41",X"49",X"08",X"09",X"01",X"12",X"6E",X"93",X"06",
		X"04",X"6E",X"EA",X"B5",X"B5",X"20",X"47",X"80",X"47",X"09",X"9F",X"08",X"41",X"93",X"10",X"6E",
		X"01",X"EA",X"04",X"6E",X"06",X"47",X"B5",X"20",X"B5",X"E0",X"47",X"09",X"80",X"11",X"41",X"93",
		X"08",X"04",X"01",X"EA",X"6E",X"B5",X"06",X"47",X"6E",X"47",X"B5",X"3E",X"20",X"41",X"80",X"10",
		X"09",X"01",X"08",X"04",X"93",X"06",X"6E",X"B5",X"EA",X"B5",X"6E",X"47",X"47",X"80",X"20",X"41",
		X"43",X"08",X"09",X"01",X"13",X"6E",X"93",X"06",X"04",X"6E",X"EA",X"B5",X"B5",X"20",X"47",X"80",
		X"47",X"09",X"52",X"08",X"41",X"93",X"11",X"6E",X"01",X"EA",X"04",X"6E",X"06",X"47",X"B5",X"40",
		X"B5",X"E3",X"47",X"09",X"80",X"10",X"41",X"97",X"08",X"27",X"01",X"EA",X"6E",X"B5",X"06",X"47",
		X"6E",X"47",X"B5",X"7D",X"20",X"41",X"80",X"10",X"09",X"01",X"08",X"41",X"D6",X"06",X"6E",X"B5",
		X"EA",X"B5",X"6E",X"47",X"47",X"4C",X"01",X"09",X"F3",X"92",X"B3",X"23",X"34",X"BE",X"3E",X"B5",
		X"73",X"B5",X"6E",X"47",X"42",X"4C",X"07",X"09",X"F3",X"92",X"B3",X"23",X"34",X"BE",X"3E",X"6E",
		X"10",X"41",X"9A",X"14",X"B5",X"10",X"46",X"09",X"D7",X"06",X"6E",X"B5",X"20",X"64",X"43",X"D0",
		X"47",X"09",X"87",X"20",X"41",X"F1",X"16",X"6E",X"24",X"D0",X"05",X"41",X"06",X"47",X"B5",X"52",
		X"14",X"6E",X"F0",X"06",X"09",X"07",X"20",X"64",X"B5",X"70",X"47",X"09",X"D0",X"14",X"41",X"F1",
		X"20",X"64",X"03",X"D0",X"6E",X"B5",X"06",X"47",X"41",X"F2",X"14",X"6E",X"73",X"20",X"09",X"03",
		X"06",X"47",X"B5",X"92",X"64",X"41",X"D0",X"10",X"09",X"01",X"08",X"43",X"F9",X"06",X"6E",X"B5",
		X"EA",X"11",X"41",X"24",X"47",X"09",X"31",X"09",X"6E",X"B5",X"06",X"47",X"20",X"EA",X"24",X"41",
		X"44",X"09",X"09",X"01",X"11",X"6E",X"3C",X"06",X"40",X"41",X"EA",X"10",X"B5",X"D6",X"47",X"09",
		X"7C",X"06",X"6E",X"B5",X"09",X"45",X"01",X"EA",X"47",X"FE",X"99",X"08",X"6A",X"01",X"34",X"27",
		X"41",X"C1",X"11",X"6E",X"61",X"09",X"09",X"01",X"06",X"47",X"B5",X"08",X"27",X"60",X"EA",X"FE",
		X"02",X"61",X"27",X"09",X"08",X"11",X"41",X"88",X"09",X"27",X"01",X"EA",X"6E",X"B5",X"06",X"47",
		X"60",X"11",X"41",X"AF",X"25",X"09",X"61",X"09",X"6E",X"B5",X"06",X"47",X"01",X"EA",X"27",X"41",
		X"E4",X"09",X"09",X"01",X"10",X"6E",X"EE",X"06",X"61",X"6A",X"EA",X"34",X"B5",X"BB",X"47",X"FE",
		X"00",X"7C",X"27",X"09",X"08",X"11",X"41",X"D7",X"09",X"06",X"01",X"EA",X"6E",X"B5",X"06",X"47",
		X"60",X"08",X"FE",X"41",X"4B",X"27",X"01",X"7C",X"11",X"6E",X"F5",X"06",X"09",X"01",X"09",X"06",
		X"B5",X"08",X"47",X"02",X"EA",X"FE",X"60",X"08",X"27",X"09",X"7C",X"09",X"41",X"9B",X"11",X"6E",
		X"01",X"EA",X"05",X"60",X"06",X"47",X"B5",X"25",X"41",X"B8",X"11",X"6E",X"7C",X"09",X"09",X"01",
		X"06",X"47",X"B5",X"92",X"05",X"6E",X"EA",X"4A",X"1E",X"4A",X"6E",X"34",X"11",X"AA",X"7C",X"6E",
		X"6B",X"6E",X"AB",X"4A",X"4A",X"44",X"34",X"AC",X"34",X"AD",X"21",X"6E",X"6E",X"34",X"4A",X"04",
		X"B5",X"4A",X"47",X"34",X"4C",X"AA",X"AF",X"09",X"F3",X"08",X"B3",X"B5",X"34",X"10",X"3E",X"F6",
		X"0B",X"B5",X"D2",X"0B",X"B5",X"9E",X"0B",X"B5",X"D6",X"0B",X"B5",X"4A",X"0B",X"AF",X"BA",X"75",
		X"35",X"4A",X"78",X"35",X"4A",X"C3",X"35",X"4A",X"AE",X"35",X"4A",X"9C",X"35",X"4A",X"B1",X"35",
		X"4A",X"FA",X"35",X"4A",X"FF",X"47",X"B5",X"90",X"50",X"B3",X"F3",X"08",X"09",X"3E",X"34",X"26",
		X"09",X"36",X"34",X"02",X"F4",X"08",X"B3",X"60",X"B6",X"8C",X"A6",X"B5",X"B3",X"07",X"93",X"BF",
		X"47",X"B3",X"F3",X"B3",X"09",X"9E",X"34",X"AE",X"09",X"A6",X"34",X"C6",X"F4",X"B3",X"B3",X"B3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"34",X"4E",X"37",X"BD",X"01",X"FF",X"00",X"C8",X"6E",X"50",X"4A",X"F5",X"FF",X"09",X"01",X"34",
		X"FF",X"08",X"9C",X"BE",X"BE",X"9C",X"08",X"FF",X"FF",X"01",X"63",X"77",X"77",X"63",X"01",X"FF",
		X"BE",X"08",X"88",X"9C",X"9C",X"88",X"08",X"BE",X"77",X"01",X"41",X"63",X"63",X"41",X"01",X"77",
		X"88",X"08",X"88",X"88",X"88",X"88",X"08",X"88",X"41",X"01",X"41",X"41",X"41",X"41",X"01",X"41",
		X"15",X"2C",X"15",X"1F",X"59",X"13",X"53",X"50",X"59",X"18",X"19",X"20",X"52",X"54",X"17",X"61",
		X"69",X"19",X"62",X"19",X"68",X"17",X"14",X"54",X"52",X"54",X"58",X"13",X"15",X"15",X"20",X"18",
		X"53",X"4A",X"11",X"34",X"54",X"98",X"52",X"6A",X"9B",X"0F",X"D6",X"9B",X"34",X"4A",X"01",X"34",
		X"09",X"9E",X"34",X"B8",X"F4",X"6A",X"B3",X"34",X"4A",X"43",X"34",X"6A",X"BC",X"00",X"B5",X"99",
		X"34",X"0C",X"00",X"B5",X"FE",X"25",X"B2",X"02",X"47",X"FE",X"0C",X"48",X"93",X"04",X"25",X"29",
		X"41",X"BD",X"11",X"6E",X"26",X"67",X"09",X"01",X"06",X"47",X"B5",X"40",X"41",X"41",X"EA",X"12",
		X"09",X"01",X"67",X"02",X"FE",X"06",X"6E",X"B5",X"EA",X"11",X"41",X"9A",X"47",X"09",X"5A",X"67",
		X"6E",X"B5",X"06",X"47",X"01",X"EA",X"23",X"60",X"C4",X"09",X"C0",X"08",X"41",X"00",X"10",X"6E",
		X"01",X"EA",X"61",X"60",X"06",X"47",X"B5",X"85",X"6A",X"5F",X"50",X"4B",X"10",X"08",X"B3",X"6A",
		X"99",X"28",X"FE",X"6A",X"34",X"45",X"00",X"98",X"34",X"0D",X"04",X"04",X"FE",X"D6",X"68",X"4A",
		X"98",X"34",X"6A",X"02",X"34",X"D6",X"9B",X"0F",X"4A",X"F4",X"34",X"B3",X"9B",X"34",X"09",X"8E",
		X"6A",X"BC",X"34",X"4A",X"B8",X"34",X"4A",X"BD",X"34",X"B5",X"43",X"00",X"B5",X"0C",X"00",X"93",
		X"A6",X"50",X"4A",X"F3",X"24",X"09",X"90",X"34",X"B3",X"93",X"08",X"24",X"5E",X"75",X"03",X"B3",
		X"CE",X"AF",X"4C",X"BE",X"93",X"09",X"24",X"34",X"41",X"05",X"34",X"5F",X"BF",X"00",X"01",X"BD",
		X"C8",X"4A",X"DD",X"34",X"4A",X"DE",X"34",X"6E",X"10",X"41",X"9C",X"13",X"09",X"9D",X"13",X"01",
		X"05",X"C8",X"5F",X"DE",X"00",X"09",X"BD",X"13",X"41",X"05",X"13",X"5F",X"DF",X"00",X"01",X"BD",
		X"C8",X"13",X"4A",X"DE",X"AF",X"4A",X"9C",X"13",X"B5",X"02",X"0B",X"09",X"9A",X"0C",X"B5",X"F5",
		X"34",X"F4",X"B6",X"B3",X"B3",X"34",X"09",X"1E",X"28",X"6E",X"60",X"4A",X"02",X"00",X"62",X"03",
		X"50",X"41",X"29",X"11",X"B5",X"50",X"47",X"09",X"61",X"06",X"6E",X"B5",X"08",X"25",X"01",X"EA",
		X"47",X"4C",X"03",X"09",X"6E",X"47",X"B5",X"F4",X"34",X"BC",X"BE",X"6D",X"B3",X"34",X"6A",X"4A",
		X"BC",X"09",X"6E",X"10",X"34",X"46",X"10",X"41",X"47",X"00",X"01",X"BD",X"10",X"5F",X"20",X"C8",
		X"B5",X"DE",X"00",X"93",X"43",X"0B",X"B5",X"0C",X"26",X"B3",X"F4",X"08",X"09",X"1E",X"34",X"D6",
		X"B3",X"6A",X"28",X"34",X"3E",X"F4",X"E8",X"B3",X"7F",X"29",X"4F",X"41",X"08",X"47",X"B5",X"50",
		X"11",X"6E",X"0E",X"06",X"09",X"01",X"08",X"25",X"B5",X"03",X"47",X"4C",X"EA",X"B5",X"6E",X"47",
		X"09",X"AE",X"34",X"BD",X"F4",X"6A",X"B3",X"34",X"6D",X"6E",X"BD",X"09",X"4A",X"10",X"34",X"02",
		X"10",X"01",X"03",X"00",X"41",X"20",X"10",X"5F",X"BD",X"00",X"B5",X"FE",X"C8",X"B5",X"0C",X"0B",
		X"60",X"4A",X"6E",X"50",X"4A",X"03",X"01",X"60",X"92",X"09",X"29",X"34",X"B5",X"F4",X"47",X"B3",
		X"1E",X"40",X"A0",X"09",X"08",X"11",X"41",X"4B",X"08",X"41",X"01",X"EA",X"6E",X"B5",X"06",X"47",
		X"09",X"96",X"35",X"01",X"75",X"6E",X"B3",X"B5",X"4C",X"34",X"09",X"3E",X"47",X"B3",X"F4",X"28",
		X"CC",X"B5",X"A3",X"0B",X"93",X"9E",X"25",X"09",X"F5",X"28",X"B3",X"B3",X"34",X"43",X"36",X"A6",
		X"09",X"96",X"35",X"90",X"FF",X"4A",X"B3",X"50",X"6A",X"00",X"35",X"DE",X"FF",X"08",X"FE",X"60",
		X"05",X"4C",X"02",X"09",X"6E",X"47",X"B5",X"9C",X"35",X"BA",X"96",X"B5",X"B3",X"0B",X"B5",X"FA",
		X"47",X"B3",X"F4",X"28",X"09",X"36",X"34",X"DB",X"B3",X"B5",X"6E",X"47",X"A6",X"4C",X"01",X"B5",
		X"BF",X"34",X"09",X"56",X"47",X"B3",X"F4",X"08",X"27",X"B5",X"BE",X"47",X"B5",X"BF",X"0B",X"09",
		X"F4",X"08",X"B3",X"60",X"34",X"21",X"76",X"67",X"B3",X"0C",X"B5",X"BA",X"C6",X"60",X"26",X"B3",
		X"E6",X"B3",X"F5",X"09",X"09",X"B6",X"34",X"F4",X"34",X"05",X"3E",X"22",X"B3",X"B5",X"08",X"0C",
		X"60",X"0C",X"B5",X"A5",X"C2",X"60",X"06",X"6A",X"DC",X"08",X"FE",X"09",X"34",X"2E",X"00",X"F4",
		X"34",X"2F",X"3E",X"BD",X"B3",X"6A",X"08",X"34",X"FE",X"B5",X"08",X"47",X"00",X"29",X"36",X"41",
		X"C0",X"08",X"09",X"01",X"11",X"6E",X"14",X"06",X"21",X"6E",X"EA",X"B5",X"B5",X"02",X"47",X"4C",
		X"47",X"09",X"D3",X"34",X"B5",X"F3",X"43",X"B3",X"DE",X"D6",X"7C",X"4A",X"93",X"01",X"07",X"DC",
		X"34",X"6A",X"F9",X"34",X"93",X"BC",X"25",X"FE",X"00",X"F4",X"0D",X"B3",X"08",X"34",X"09",X"1E",
		X"08",X"47",X"B5",X"D8",X"B2",X"41",X"29",X"10",X"09",X"01",X"08",X"44",X"35",X"06",X"6E",X"B5",
		X"EA",X"B5",X"6E",X"47",X"47",X"4C",X"03",X"93",X"CC",X"0B",X"B5",X"A9",X"25",X"93",X"FA",X"25",
		X"B5",X"A9",X"0B",X"2A",X"DA",X"25",X"93",X"D7",X"34",X"00",X"F5",X"F5",X"BB",X"00",X"09",X"61",
		X"F5",X"86",X"01",X"17",X"7E",X"02",X"F5",X"9E",X"27",X"B3",X"5F",X"B3",X"F5",X"68",X"02",X"68",
		X"B3",X"F5",X"B3",X"00",X"68",X"7E",X"68",X"09",X"4C",X"B5",X"B3",X"47",X"27",X"C5",X"0F",X"76",
		X"0B",X"10",X"BB",X"10",X"56",X"27",X"B9",X"27",X"11",X"51",X"31",X"71",X"27",X"27",X"27",X"27",
		X"B1",X"C0",X"7E",X"5F",X"F5",X"F5",X"04",X"04",X"B1",X"80",X"7E",X"5F",X"F5",X"F5",X"04",X"04",
		X"B1",X"80",X"7E",X"5F",X"F5",X"F5",X"03",X"03",X"B1",X"C0",X"7E",X"5F",X"F5",X"F5",X"03",X"03",
		X"B1",X"BB",X"8C",X"09",X"2A",X"F5",X"34",X"00",X"00",X"01",X"61",X"34",X"F5",X"00",X"BB",X"4F",
		X"6F",X"F5",X"12",X"00",X"BD",X"7E",X"9D",X"09",X"84",X"B5",X"B3",X"47",X"27",X"C5",X"0F",X"76",
		X"0B",X"54",X"BB",X"C0",X"56",X"40",X"B9",X"27",X"D3",X"3D",X"1B",X"80",X"27",X"40",X"40",X"40",
		X"F5",X"8A",X"03",X"F5",X"7E",X"34",X"4A",X"7E",X"04",X"B5",X"8B",X"40",X"4A",X"BA",X"34",X"F5",
		X"7E",X"50",X"42",X"FE",X"06",X"34",X"6A",X"00",X"08",X"34",X"6A",X"00",X"47",X"FE",X"51",X"08",
		X"47",X"34",X"09",X"9D",X"91",X"21",X"52",X"D1",X"43",X"4E",X"05",X"BD",X"01",X"FF",X"00",X"C8",
		X"B1",X"43",X"7E",X"60",X"F5",X"42",X"06",X"B9",X"F5",X"08",X"06",X"61",X"7E",X"00",X"09",X"BB",
		X"42",X"42",X"F6",X"F5",X"60",X"41",X"B5",X"7E",X"03",X"34",X"4A",X"7E",X"C0",X"F5",X"8A",X"04",
		X"4A",X"BA",X"34",X"6A",X"8B",X"40",X"B5",X"50",X"34",X"4A",X"00",X"50",X"FE",X"6A",X"28",X"34",
		X"B3",X"05",X"F5",X"6D",X"0F",X"80",X"16",X"91",X"FD",X"FD",X"52",X"FD",X"09",X"21",X"34",X"5B",
		X"CC",X"EE",X"11",X"11",X"33",X"EE",X"CC",X"00",X"11",X"33",X"66",X"44",X"44",X"33",X"11",X"00",
		X"11",X"11",X"FF",X"FF",X"11",X"11",X"00",X"00",X"00",X"00",X"77",X"77",X"22",X"00",X"00",X"00",
		X"11",X"99",X"DD",X"DD",X"FF",X"77",X"33",X"00",X"33",X"77",X"55",X"44",X"44",X"66",X"22",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"33",X"22",X"00",X"44",X"66",X"77",X"55",X"44",X"44",X"00",X"00",
		X"00",X"92",X"08",X"B1",X"00",X"92",X"84",X"B1",X"00",X"64",X"01",X"78",X"00",X"64",X"42",X"78",
		X"03",X"C1",X"B2",X"9C",X"6C",X"80",X"D1",X"BE",X"0C",X"C8",X"74",X"63",X"93",X"40",X"E8",X"77",
		X"B1",X"84",X"92",X"00",X"B1",X"08",X"92",X"00",X"78",X"42",X"64",X"00",X"78",X"01",X"64",X"00",
		X"FF",X"F1",X"F7",X"6C",X"F7",X"F0",X"F3",X"03",X"FF",X"F8",X"FE",X"93",X"FE",X"F0",X"FC",X"0C",
		X"00",X"92",X"08",X"B1",X"00",X"92",X"84",X"B1",X"00",X"25",X"01",X"39",X"00",X"25",X"42",X"39",
		X"03",X"63",X"F3",X"00",X"6C",X"41",X"FF",X"36",X"0C",X"FE",X"F8",X"FF",X"93",X"FF",X"FC",X"FF",
		X"B1",X"84",X"92",X"00",X"B1",X"08",X"92",X"00",X"39",X"42",X"25",X"00",X"39",X"01",X"25",X"00",
		X"36",X"FF",X"41",X"6C",X"00",X"F3",X"63",X"03",X"FF",X"FC",X"FF",X"93",X"FF",X"F8",X"FE",X"0C",
		X"00",X"9A",X"08",X"21",X"00",X"16",X"84",X"A9",X"00",X"64",X"01",X"78",X"00",X"64",X"42",X"78",
		X"03",X"93",X"F0",X"0F",X"6C",X"87",X"93",X"0F",X"0C",X"0C",X"6C",X"00",X"93",X"08",X"6F",X"41",
		X"A9",X"84",X"16",X"00",X"21",X"08",X"9A",X"00",X"78",X"42",X"64",X"00",X"78",X"01",X"64",X"00",
		X"0F",X"93",X"87",X"6C",X"0F",X"F0",X"93",X"03",X"41",X"6F",X"08",X"93",X"00",X"6C",X"0C",X"0C",
		X"00",X"92",X"08",X"B1",X"00",X"92",X"84",X"B1",X"00",X"64",X"01",X"78",X"00",X"64",X"42",X"78",
		X"03",X"0F",X"93",X"0F",X"6C",X"0F",X"0F",X"0F",X"0C",X"8E",X"78",X"0F",X"93",X"8E",X"6C",X"0F",
		X"B1",X"84",X"92",X"00",X"B1",X"08",X"92",X"00",X"78",X"42",X"64",X"00",X"78",X"01",X"64",X"00",
		X"0F",X"0F",X"0F",X"6C",X"0F",X"93",X"0F",X"03",X"0F",X"6C",X"8E",X"93",X"0F",X"78",X"8E",X"0C",
		X"00",X"92",X"08",X"B1",X"00",X"92",X"84",X"B1",X"00",X"64",X"01",X"78",X"00",X"64",X"42",X"78",
		X"03",X"B6",X"F0",X"88",X"6C",X"94",X"F3",X"C9",X"0C",X"76",X"F0",X"41",X"93",X"62",X"FC",X"C9",
		X"B1",X"84",X"92",X"00",X"B1",X"08",X"92",X"00",X"78",X"42",X"64",X"00",X"78",X"01",X"64",X"00",
		X"C9",X"F3",X"94",X"6C",X"88",X"F0",X"B6",X"03",X"C9",X"FC",X"62",X"93",X"41",X"F0",X"76",X"0C",
		X"00",X"B0",X"80",X"F0",X"00",X"B0",X"90",X"F0",X"00",X"02",X"01",X"0A",X"00",X"06",X"00",X"0A",
		X"43",X"49",X"2C",X"0C",X"4E",X"0C",X"59",X"06",X"90",X"C8",X"70",X"63",X"F0",X"40",X"E8",X"77",
		X"F0",X"90",X"B0",X"00",X"F0",X"80",X"B0",X"00",X"0B",X"0B",X"0D",X"03",X"05",X"07",X"0B",X"00",
		X"47",X"0D",X"0B",X"01",X"03",X"0B",X"09",X"00",X"FF",X"78",X"FE",X"6C",X"FE",X"6C",X"7C",X"18",
		X"00",X"B0",X"80",X"FC",X"00",X"B8",X"90",X"FC",X"00",X"03",X"00",X"0F",X"00",X"07",X"00",X"07",
		X"00",X"0C",X"03",X"00",X"01",X"08",X"4F",X"36",X"08",X"FF",X"FC",X"63",X"78",X"77",X"FE",X"63",
		X"FC",X"90",X"B8",X"00",X"FC",X"80",X"B0",X"00",X"0D",X"00",X"07",X"00",X"0F",X"00",X"03",X"00",
		X"36",X"4F",X"08",X"01",X"00",X"03",X"0C",X"00",X"63",X"FE",X"77",X"78",X"63",X"FC",X"FF",X"08",
		X"00",X"B8",X"80",X"60",X"00",X"34",X"90",X"E8",X"00",X"03",X"00",X"0E",X"00",X"07",X"00",X"07",
		X"00",X"0D",X"03",X"4F",X"01",X"03",X"0E",X"4F",X"0C",X"9C",X"7C",X"00",X"78",X"88",X"FF",X"41",
		X"E8",X"90",X"34",X"00",X"60",X"80",X"B8",X"00",X"0D",X"00",X"07",X"00",X"0E",X"00",X"03",X"00",
		X"4F",X"0F",X"03",X"01",X"4F",X"03",X"0D",X"00",X"41",X"FF",X"88",X"78",X"00",X"7C",X"9C",X"0C",
		X"00",X"B0",X"80",X"F8",X"00",X"B8",X"90",X"F8",X"00",X"03",X"00",X"0E",X"00",X"07",X"01",X"0F",
		X"01",X"0E",X"47",X"0C",X"03",X"0C",X"4F",X"4D",X"90",X"77",X"FC",X"41",X"F0",X"63",X"FE",X"C9",
		X"F8",X"90",X"B8",X"00",X"F8",X"80",X"B0",X"00",X"0D",X"01",X"07",X"00",X"0E",X"00",X"03",X"00",
		X"4D",X"4F",X"0C",X"03",X"0C",X"47",X"0E",X"01",X"C9",X"FE",X"63",X"F0",X"41",X"FC",X"77",X"90",
		X"15",X"2C",X"15",X"1F",X"59",X"13",X"53",X"50",X"59",X"18",X"19",X"20",X"52",X"54",X"17",X"61",
		X"69",X"19",X"62",X"19",X"68",X"17",X"14",X"54",X"52",X"54",X"58",X"13",X"15",X"15",X"20",X"18",
		X"53",X"84",X"11",X"EF",X"54",X"C2",X"52",X"08",X"01",X"12",X"34",X"7F",X"7F",X"34",X"12",X"01",
		X"0C",X"C2",X"E1",X"E9",X"E9",X"E1",X"C2",X"0C",X"03",X"34",X"78",X"79",X"79",X"78",X"34",X"03",
		X"0C",X"C2",X"ED",X"E5",X"E5",X"ED",X"C2",X"0C",X"03",X"34",X"7B",X"7A",X"7A",X"7B",X"34",X"03",
		X"0C",X"CE",X"E3",X"E3",X"E3",X"E3",X"CE",X"0C",X"03",X"37",X"7C",X"7C",X"7C",X"7C",X"37",X"03",
		X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"88",X"CC",X"22",X"22",X"66",X"CC",X"88",X"00",X"33",X"77",X"CC",X"88",X"88",X"77",X"33",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"00",X"00",X"FF",X"FF",X"44",X"00",X"00",X"00",
		X"22",X"22",X"AA",X"AA",X"EE",X"EE",X"66",X"00",X"66",X"FF",X"BB",X"99",X"99",X"CC",X"44",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"88",X"DD",X"FF",X"BB",X"99",X"88",X"00",X"00",
		X"88",X"EE",X"EE",X"88",X"88",X"88",X"88",X"00",X"00",X"FF",X"FF",X"CC",X"66",X"33",X"11",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"11",X"BB",X"AA",X"AA",X"AA",X"EE",X"EE",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"00",X"99",X"99",X"99",X"DD",X"77",X"33",X"00",
		X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"CC",X"EE",X"BB",X"99",X"88",X"CC",X"CC",X"00",
		X"CC",X"EE",X"AA",X"AA",X"22",X"22",X"CC",X"00",X"00",X"66",X"99",X"99",X"BB",X"FF",X"66",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"22",X"00",X"00",X"77",X"FF",X"99",X"99",X"99",X"FF",X"66",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"88",X"88",X"88",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"CC",X"77",X"33",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"EE",X"00",X"66",X"FF",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"44",X"66",X"22",X"22",X"66",X"CC",X"88",X"00",X"44",X"CC",X"88",X"88",X"CC",X"77",X"33",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"88",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"88",X"99",X"99",X"99",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"88",X"99",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"EE",X"EE",X"22",X"22",X"66",X"CC",X"88",X"00",X"99",X"99",X"99",X"88",X"CC",X"77",X"33",X"00",
		X"EE",X"EE",X"00",X"00",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"11",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"88",X"CC",X"66",X"33",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"EE",X"EE",X"00",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"77",X"33",X"77",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"77",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"00",X"88",X"88",X"88",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"FF",X"00",
		X"AA",X"CC",X"EE",X"AA",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"99",X"88",X"88",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"00",X"55",X"DD",X"99",X"99",X"FF",X"66",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"88",X"CC",X"EE",X"CC",X"88",X"00",X"00",X"FF",X"FF",X"11",X"00",X"11",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"11",X"FF",X"FF",X"00",
		X"66",X"EE",X"CC",X"88",X"CC",X"EE",X"66",X"00",X"CC",X"EE",X"77",X"33",X"77",X"EE",X"CC",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"EE",X"FF",X"11",X"11",X"FF",X"EE",X"00",X"00",
		X"22",X"22",X"22",X"AA",X"EE",X"EE",X"66",X"00",X"CC",X"EE",X"FF",X"BB",X"99",X"88",X"88",X"00",
		X"ED",X"98",X"1A",X"C0",X"50",X"09",X"48",X"50",X"11",X"49",X"50",X"01",X"27",X"00",X"1E",X"00",
		X"ED",X"98",X"1A",X"C0",X"50",X"09",X"D8",X"67",X"11",X"D9",X"67",X"01",X"27",X"00",X"1E",X"00",
		X"ED",X"98",X"1A",X"C0",X"50",X"09",X"40",X"50",X"11",X"41",X"50",X"01",X"37",X"00",X"1E",X"00",
		X"ED",X"98",X"09",X"52",X"64",X"11",X"53",X"64",X"01",X"67",X"00",X"1E",X"FF",X"ED",X"98",X"09",
		X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",
		X"CC",X"22",X"01",X"4C",X"22",X"11",X"22",X"CC",X"33",X"44",X"88",X"44",X"23",X"08",X"44",X"33",
		X"1C",X"0B",X"E5",X"95",X"17",X"7E",X"1A",X"E8",X"64",X"78",X"CE",X"18",X"09",X"DC",X"0A",X"E5",
		X"95",X"17",X"0A",X"E9",X"64",X"78",X"CE",X"18",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",X"E3",X"3F",
		X"CE",X"00",X"33",X"04",X"02",X"C0",X"00",X"37",X"00",X"11",X"22",X"22",X"22",X"33",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"44",X"44",X"44",X"88",X"00",
		X"40",X"ED",X"98",X"09",X"C2",X"47",X"11",X"C3",X"47",X"01",X"34",X"00",X"1E",X"01",X"ED",X"98",
		X"1A",X"C0",X"50",X"09",X"CA",X"47",X"11",X"CB",X"47",X"01",X"34",X"00",X"1E",X"05",X"ED",X"98",
		X"02",X"44",X"99",X"89",X"88",X"88",X"55",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"AA",X"11",X"11",X"89",X"99",X"22",X"04",
		X"00",X"ED",X"98",X"09",X"FC",X"64",X"11",X"DA",X"43",X"E5",X"05",X"12",X"09",X"02",X"40",X"11",
		X"03",X"40",X"01",X"3C",X"00",X"1E",X"40",X"ED",X"98",X"1A",X"C0",X"50",X"09",X"02",X"44",X"11",
		X"00",X"00",X"00",X"02",X"22",X"22",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"88",X"44",X"44",X"04",X"00",X"00",X"00",X"FF",X"88",X"88",X"8A",X"86",X"11",X"11",X"FF",
		X"06",X"00",X"ED",X"98",X"AF",X"1A",X"24",X"40",X"3A",X"C9",X"64",X"FE",X"00",X"08",X"23",X"09",
		X"F1",X"37",X"11",X"24",X"40",X"01",X"21",X"00",X"ED",X"98",X"1A",X"C0",X"50",X"09",X"42",X"65",
		X"11",X"43",X"65",X"01",X"FF",X"00",X"1E",X"00",X"ED",X"98",X"09",X"5B",X"32",X"0A",X"73",X"65",
		X"0A",X"43",X"65",X"09",X"72",X"65",X"0A",X"62",X"65",X"09",X"8D",X"32",X"0A",X"5E",X"65",X"0A",
		X"76",X"65",X"09",X"5D",X"65",X"0A",X"4D",X"65",X"09",X"D7",X"32",X"0A",X"91",X"65",X"0A",X"79",
		X"65",X"09",X"90",X"65",X"0A",X"80",X"65",X"09",X"21",X"33",X"0A",X"AC",X"65",X"0A",X"94",X"65",
		X"00",X"00",X"4C",X"00",X"FF",X"11",X"89",X"11",X"00",X"00",X"33",X"44",X"88",X"89",X"88",X"FF",
		X"22",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"65",X"0A",X"D1",X"65",X"09",X"B7",X"33",X"0A",X"FD",X"65",X"0A",X"CD",X"65",X"09",X"FC",X"65",
		X"0A",X"EC",X"65",X"09",X"D1",X"33",X"0A",X"30",X"66",X"0A",X"00",X"66",X"09",X"17",X"66",X"0A",
		X"00",X"00",X"00",X"00",X"44",X"AA",X"11",X"11",X"00",X"00",X"00",X"00",X"02",X"44",X"99",X"89",
		X"19",X"99",X"22",X"04",X"00",X"00",X"00",X"00",X"88",X"88",X"55",X"22",X"00",X"00",X"00",X"00",
		X"64",X"FE",X"00",X"C2",X"EE",X"23",X"09",X"F3",X"64",X"E3",X"8E",X"AF",X"1A",X"01",X"50",X"09",
		X"F4",X"64",X"E3",X"86",X"E5",X"EF",X"17",X"1A",X"C0",X"50",X"3E",X"40",X"E5",X"CA",X"16",X"3E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"22",
		X"11",X"19",X"45",X"44",X"44",X"CC",X"00",X"00",X"22",X"2A",X"81",X"88",X"44",X"33",X"00",X"00",
		X"E5",X"D0",X"17",X"11",X"35",X"47",X"09",X"E6",X"20",X"3E",X"01",X"06",X"04",X"E5",X"D0",X"17",
		X"11",X"A2",X"44",X"09",X"E7",X"20",X"3E",X"01",X"06",X"04",X"E5",X"D0",X"17",X"11",X"0E",X"46",
		X"09",X"D4",X"20",X"3E",X"01",X"06",X"04",X"E5",X"D0",X"17",X"11",X"CF",X"44",X"09",X"D6",X"20",
		X"3E",X"01",X"06",X"04",X"E5",X"D0",X"17",X"11",X"A9",X"46",X"09",X"D1",X"20",X"3E",X"01",X"06",
		X"04",X"E5",X"D0",X"17",X"11",X"A3",X"45",X"09",X"D0",X"20",X"3E",X"01",X"06",X"04",X"E5",X"D0",
		X"17",X"11",X"64",X"47",X"09",X"D5",X"20",X"3E",X"01",X"06",X"04",X"E5",X"D0",X"17",X"11",X"25",
		X"46",X"09",X"E6",X"20",X"3E",X"01",X"06",X"04",X"E5",X"D0",X"17",X"11",X"6E",X"44",X"09",X"D6",
		X"20",X"3E",X"01",X"06",X"04",X"E5",X"D0",X"17",X"11",X"E7",X"46",X"09",X"D3",X"20",X"3E",X"01",
		X"06",X"04",X"E5",X"D0",X"17",X"11",X"67",X"45",X"09",X"D2",X"20",X"3E",X"01",X"06",X"04",X"E5",
		X"D0",X"17",X"11",X"19",X"46",X"09",X"E5",X"20",X"3E",X"01",X"06",X"04",X"E5",X"D0",X"17",X"11",
		X"52",X"45",X"09",X"E6",X"20",X"3E",X"01",X"06",X"04",X"E5",X"D0",X"17",X"11",X"13",X"47",X"09",
		X"D4",X"20",X"3E",X"01",X"06",X"04",X"E5",X"D0",X"17",X"11",X"D4",X"44",X"09",X"D2",X"20",X"3E",
		X"01",X"06",X"04",X"E5",X"D0",X"17",X"11",X"15",X"46",X"09",X"E5",X"20",X"3E",X"01",X"06",X"04",
		X"E5",X"D0",X"17",X"11",X"B8",X"46",X"09",X"D3",X"20",X"3E",X"01",X"06",X"04",X"E5",X"D0",X"17",
		X"11",X"B0",X"45",X"09",X"D5",X"20",X"3E",X"01",X"06",X"04",X"E5",X"D0",X"17",X"11",X"72",X"47",
		X"09",X"E7",X"20",X"3E",X"01",X"06",X"04",X"E5",X"D0",X"17",X"C3",X"F3",X"20",X"01",X"03",X"05",
		X"07",X"21",X"26",X"27",X"10",X"30",X"36",X"12",X"03",X"05",X"07",X"11",X"67",X"41",X"09",X"C3",
		X"08",X"3E",X"01",X"06",X"04",X"E5",X"BA",X"17",X"3E",X"20",X"E5",X"80",X"17",X"11",X"0E",X"42",
		X"09",X"C3",X"08",X"3E",X"01",X"06",X"04",X"E5",X"BA",X"17",X"3E",X"20",X"E5",X"80",X"17",X"11",
		X"E7",X"42",X"09",X"C3",X"08",X"3E",X"01",X"06",X"04",X"E5",X"BA",X"17",X"3E",X"20",X"E5",X"80",
		X"17",X"11",X"A2",X"40",X"09",X"C3",X"08",X"3E",X"01",X"06",X"04",X"E5",X"BA",X"17",X"3E",X"20",
		X"E5",X"80",X"17",X"11",X"15",X"42",X"09",X"C3",X"08",X"3E",X"01",X"06",X"04",X"E5",X"BA",X"17",
		X"3E",X"20",X"E5",X"80",X"17",X"11",X"35",X"43",X"09",X"C3",X"08",X"3E",X"01",X"06",X"04",X"E5",
		X"BA",X"17",X"3E",X"20",X"E5",X"80",X"17",X"11",X"D4",X"40",X"09",X"C3",X"08",X"3E",X"01",X"06",
		X"04",X"E5",X"BA",X"17",X"3E",X"20",X"E5",X"80",X"17",X"11",X"A9",X"42",X"09",X"C3",X"08",X"3E",
		X"01",X"06",X"04",X"E5",X"BA",X"17",X"3E",X"20",X"E5",X"80",X"17",X"11",X"72",X"43",X"09",X"C3",
		X"08",X"3E",X"01",X"06",X"04",X"E5",X"BA",X"17",X"3E",X"20",X"E5",X"80",X"17",X"11",X"5F",X"40",
		X"09",X"C3",X"08",X"3E",X"01",X"06",X"04",X"E5",X"BA",X"17",X"3E",X"20",X"E5",X"80",X"17",X"11",
		X"A3",X"41",X"09",X"C3",X"08",X"3E",X"01",X"06",X"04",X"E5",X"BA",X"17",X"3E",X"20",X"E5",X"80",
		X"17",X"11",X"64",X"43",X"09",X"C3",X"08",X"3E",X"01",X"06",X"04",X"E5",X"BA",X"17",X"3E",X"20",
		X"E5",X"80",X"17",X"11",X"25",X"42",X"09",X"C3",X"08",X"3E",X"01",X"06",X"04",X"E5",X"BA",X"17",
		X"3E",X"20",X"E5",X"80",X"17",X"11",X"B8",X"42",X"09",X"C3",X"08",X"3E",X"01",X"06",X"04",X"E5",
		X"BA",X"17",X"3E",X"20",X"E5",X"80",X"17",X"11",X"19",X"42",X"09",X"C3",X"08",X"3E",X"01",X"06",
		X"04",X"E5",X"BA",X"17",X"3E",X"20",X"E5",X"80",X"17",X"11",X"CF",X"40",X"09",X"C3",X"08",X"3E",
		X"01",X"06",X"04",X"E5",X"BA",X"17",X"3E",X"20",X"E5",X"80",X"17",X"11",X"B0",X"41",X"09",X"C3",
		X"08",X"3E",X"01",X"06",X"04",X"E5",X"BA",X"17",X"3E",X"20",X"E5",X"80",X"17",X"11",X"6E",X"40",
		X"09",X"C3",X"08",X"3E",X"01",X"06",X"04",X"E5",X"BA",X"17",X"3E",X"20",X"E5",X"80",X"17",X"11",
		X"13",X"43",X"09",X"C3",X"08",X"3E",X"01",X"06",X"04",X"E5",X"BA",X"17",X"3E",X"20",X"E5",X"80",
		X"17",X"11",X"52",X"41",X"09",X"C3",X"08",X"3E",X"01",X"06",X"04",X"E5",X"BA",X"17",X"3E",X"10",
		X"E5",X"80",X"17",X"11",X"B3",X"40",X"09",X"C7",X"08",X"3E",X"01",X"06",X"27",X"E5",X"BA",X"17",
		X"3E",X"20",X"E5",X"80",X"17",X"11",X"7D",X"40",X"09",X"D6",X"08",X"3E",X"01",X"06",X"11",X"E5",
		X"BA",X"17",X"3E",X"01",X"E5",X"1C",X"17",X"09",X"F3",X"64",X"E3",X"6E",X"C2",X"EE",X"23",X"E5",
		X"73",X"12",X"3E",X"07",X"E5",X"1C",X"17",X"09",X"F3",X"64",X"E3",X"6E",X"C2",X"EE",X"23",X"3E",
		X"40",X"E5",X"CA",X"16",X"11",X"40",X"44",X"09",X"D7",X"20",X"3E",X"13",X"06",X"34",X"E5",X"D0",
		X"17",X"11",X"87",X"46",X"09",X"F1",X"20",X"3E",X"24",X"06",X"05",X"E5",X"D0",X"17",X"11",X"52",
		X"44",X"09",X"F0",X"20",X"3E",X"07",X"06",X"34",X"E5",X"D0",X"17",X"11",X"70",X"44",X"09",X"F1",
		X"20",X"3E",X"03",X"06",X"34",X"E5",X"D0",X"17",X"11",X"73",X"44",X"09",X"F2",X"20",X"3E",X"03",
		X"06",X"34",X"E5",X"D0",X"17",X"11",X"C2",X"40",X"09",X"F9",X"08",X"3E",X"01",X"06",X"13",X"E5",
		X"BA",X"17",X"11",X"61",X"41",X"09",X"24",X"09",X"3E",X"20",X"06",X"24",X"E5",X"BA",X"17",X"11",
		X"14",X"41",X"09",X"6C",X"09",X"3E",X"01",X"06",X"10",X"E5",X"BA",X"17",X"11",X"D6",X"40",X"09",
		X"7C",X"09",X"3E",X"01",X"06",X"15",X"E5",X"BA",X"17",X"3A",X"C9",X"64",X"FE",X"01",X"08",X"27",
		X"11",X"31",X"41",X"09",X"91",X"09",X"3E",X"01",X"06",X"27",X"E5",X"BA",X"17",X"30",X"08",X"FE",
		X"02",X"08",X"27",X"11",X"31",X"41",X"09",X"88",X"09",X"3E",X"01",X"06",X"27",X"E5",X"BA",X"17",
		X"30",X"25",X"11",X"31",X"41",X"09",X"AF",X"09",X"3E",X"01",X"06",X"27",X"E5",X"BA",X"17",X"11",
		X"B4",X"40",X"09",X"BE",X"09",X"3E",X"01",X"06",X"31",X"E5",X"BA",X"17",X"3A",X"EB",X"64",X"FE",
		X"00",X"08",X"27",X"11",X"7C",X"41",X"09",X"D7",X"09",X"3E",X"01",X"06",X"06",X"E5",X"BA",X"17",
		X"30",X"1B",X"FE",X"01",X"08",X"27",X"11",X"7C",X"41",X"09",X"F5",X"09",X"3E",X"01",X"06",X"06",
		X"E5",X"BA",X"17",X"30",X"08",X"FE",X"02",X"08",X"27",X"11",X"7C",X"41",X"09",X"CB",X"09",X"3E",
		X"01",X"06",X"05",X"E5",X"BA",X"17",X"30",X"25",X"11",X"7C",X"41",X"09",X"E8",X"09",X"3E",X"01",
		X"06",X"05",X"E5",X"BA",X"17",X"3E",X"C2",X"1A",X"4E",X"41",X"3E",X"7C",X"1A",X"AA",X"64",X"3E",
		X"3B",X"1A",X"AB",X"64",X"3E",X"14",X"1A",X"AC",X"64",X"3E",X"21",X"1A",X"AD",X"64",X"3E",X"04",
		X"E5",X"1C",X"17",X"AF",X"1A",X"AA",X"64",X"09",X"F3",X"64",X"E3",X"6E",X"08",X"40",X"E5",X"F6",
		X"0B",X"E5",X"D2",X"0B",X"E5",X"CE",X"0B",X"E5",X"D6",X"0B",X"E5",X"EA",X"0B",X"AF",X"1A",X"75",
		X"65",X"1A",X"78",X"65",X"1A",X"93",X"65",X"1A",X"AE",X"65",X"1A",X"E1",X"65",X"1A",X"CC",X"65",
		X"1A",X"FF",X"65",X"E5",X"FA",X"17",X"1A",X"C0",X"50",X"09",X"F3",X"64",X"E3",X"6E",X"08",X"26",
		X"09",X"F4",X"64",X"E3",X"66",X"08",X"02",X"30",X"E6",X"E3",X"A6",X"C3",X"8C",X"07",X"E5",X"EF",
		X"17",X"09",X"F3",X"64",X"E3",X"CE",X"E3",X"AE",X"09",X"F4",X"64",X"E3",X"A6",X"E3",X"96",X"E3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"64",X"01",X"67",X"00",X"1E",X"FF",X"ED",X"98",X"3E",X"FF",X"1A",X"01",X"50",X"09",X"F5",X"64",
		X"FF",X"EE",X"CC",X"08",X"08",X"CC",X"EE",X"FF",X"FF",X"77",X"33",X"01",X"01",X"33",X"77",X"FF",
		X"EE",X"CC",X"88",X"08",X"08",X"88",X"CC",X"EE",X"77",X"33",X"11",X"01",X"01",X"11",X"33",X"77",
		X"88",X"88",X"88",X"08",X"08",X"88",X"88",X"88",X"11",X"11",X"11",X"01",X"01",X"11",X"11",X"11",
		X"45",X"59",X"45",X"53",X"2C",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",
		X"39",X"38",X"32",X"44",X"49",X"47",X"49",X"54",X"52",X"45",X"58",X"20",X"54",X"45",X"43",X"48",
		X"53",X"54",X"41",X"52",X"1A",X"C8",X"64",X"3A",X"CB",X"64",X"D6",X"01",X"0F",X"1A",X"CB",X"64",
		X"09",X"F4",X"64",X"E3",X"CE",X"3A",X"E8",X"64",X"1A",X"EC",X"64",X"E5",X"13",X"00",X"3A",X"C9",
		X"64",X"FE",X"00",X"E2",X"0C",X"25",X"E5",X"02",X"17",X"C3",X"0C",X"25",X"FE",X"04",X"18",X"29",
		X"11",X"26",X"41",X"09",X"ED",X"37",X"3E",X"01",X"06",X"11",X"E5",X"BA",X"17",X"11",X"10",X"42",
		X"09",X"FE",X"37",X"3E",X"01",X"06",X"02",X"E5",X"BA",X"17",X"11",X"5A",X"41",X"09",X"CA",X"37",
		X"3E",X"01",X"06",X"23",X"E5",X"BA",X"17",X"30",X"94",X"11",X"90",X"40",X"09",X"00",X"08",X"3E",
		X"01",X"06",X"31",X"E5",X"BA",X"17",X"30",X"85",X"3A",X"40",X"50",X"E3",X"5F",X"08",X"1B",X"3A",
		X"C9",X"64",X"FE",X"00",X"28",X"15",X"3A",X"C8",X"64",X"FE",X"04",X"38",X"0D",X"D6",X"04",X"1A",
		X"C8",X"64",X"3A",X"CB",X"64",X"D6",X"02",X"0F",X"1A",X"CB",X"64",X"09",X"F4",X"64",X"E3",X"8E",
		X"3A",X"E8",X"64",X"1A",X"EC",X"64",X"1A",X"ED",X"64",X"E5",X"13",X"00",X"E5",X"0C",X"00",X"C3",
		X"A6",X"24",X"1A",X"C0",X"50",X"09",X"F3",X"64",X"E3",X"5E",X"08",X"03",X"C3",X"75",X"24",X"E3",
		X"9E",X"C3",X"1C",X"24",X"AF",X"09",X"EE",X"64",X"11",X"EF",X"64",X"01",X"05",X"00",X"5F",X"ED",
		X"98",X"1A",X"DD",X"64",X"1A",X"DE",X"64",X"3E",X"40",X"09",X"CC",X"43",X"11",X"CD",X"43",X"01",
		X"05",X"00",X"5F",X"ED",X"98",X"09",X"DE",X"43",X"11",X"DF",X"43",X"01",X"05",X"00",X"5F",X"ED",
		X"98",X"AF",X"1A",X"CC",X"43",X"1A",X"DE",X"43",X"E5",X"CA",X"0B",X"E5",X"02",X"0C",X"09",X"F5",
		X"64",X"E3",X"E6",X"09",X"F4",X"64",X"E3",X"4E",X"28",X"02",X"30",X"32",X"3E",X"00",X"1A",X"03",
		X"50",X"E5",X"29",X"17",X"11",X"50",X"41",X"09",X"31",X"08",X"3E",X"01",X"06",X"25",X"E5",X"BA",
		X"17",X"3E",X"03",X"E5",X"1C",X"17",X"09",X"F4",X"64",X"E3",X"EE",X"3A",X"EC",X"64",X"3D",X"1A",
		X"EC",X"64",X"3E",X"40",X"09",X"16",X"40",X"11",X"17",X"40",X"01",X"20",X"00",X"5F",X"ED",X"98",
		X"E5",X"13",X"00",X"E5",X"DE",X"0B",X"C3",X"0C",X"26",X"09",X"F4",X"64",X"E3",X"4E",X"08",X"D6",
		X"E3",X"6E",X"28",X"B8",X"3A",X"F4",X"64",X"E3",X"7F",X"08",X"1F",X"E5",X"29",X"17",X"11",X"50",
		X"41",X"09",X"0E",X"08",X"3E",X"01",X"06",X"25",X"E5",X"BA",X"17",X"3E",X"03",X"E5",X"1C",X"17",
		X"09",X"F4",X"64",X"E3",X"AE",X"3A",X"ED",X"64",X"3D",X"1A",X"ED",X"64",X"3E",X"40",X"09",X"02",
		X"40",X"11",X"03",X"40",X"01",X"20",X"00",X"5F",X"ED",X"98",X"E5",X"0C",X"00",X"E5",X"FE",X"0B",
		X"30",X"1A",X"3E",X"01",X"1A",X"03",X"50",X"30",X"C2",X"E5",X"29",X"17",X"09",X"F4",X"64",X"E3",
		X"4E",X"08",X"A0",X"11",X"10",X"41",X"09",X"1B",X"08",X"3E",X"01",X"06",X"11",X"E5",X"BA",X"17",
		X"09",X"75",X"65",X"E3",X"C6",X"3E",X"01",X"E5",X"1C",X"17",X"09",X"F4",X"64",X"E3",X"6E",X"28",
		X"9C",X"C3",X"A3",X"25",X"E5",X"CE",X"0B",X"09",X"F5",X"64",X"E3",X"66",X"28",X"13",X"E3",X"A6",
		X"09",X"FF",X"65",X"E3",X"C6",X"1A",X"C0",X"50",X"3A",X"FF",X"65",X"FE",X"00",X"08",X"DE",X"30",
		X"05",X"3E",X"02",X"E5",X"1C",X"17",X"09",X"CC",X"65",X"E3",X"C6",X"E5",X"EA",X"0B",X"E5",X"FA",
		X"17",X"09",X"F4",X"64",X"E3",X"66",X"28",X"DB",X"E3",X"A6",X"3E",X"01",X"E5",X"1C",X"17",X"E5",
		X"EF",X"17",X"09",X"F4",X"64",X"E3",X"56",X"08",X"27",X"E5",X"EE",X"0B",X"E5",X"EF",X"17",X"09",
		X"F4",X"64",X"E3",X"76",X"08",X"21",X"30",X"37",X"E3",X"96",X"E5",X"26",X"0C",X"30",X"EA",X"E3",
		X"B6",X"09",X"F5",X"64",X"E3",X"E6",X"09",X"F4",X"64",X"E3",X"6E",X"08",X"05",X"E5",X"22",X"0C",
		X"30",X"92",X"E5",X"06",X"0C",X"30",X"A5",X"3A",X"DC",X"64",X"FE",X"00",X"08",X"2E",X"09",X"F4",
		X"64",X"E3",X"6E",X"08",X"2F",X"3A",X"ED",X"64",X"FE",X"00",X"08",X"66",X"E5",X"29",X"17",X"11",
		X"90",X"41",X"09",X"44",X"08",X"3E",X"01",X"06",X"21",X"E5",X"BA",X"17",X"3E",X"02",X"E5",X"1C",
		X"17",X"E5",X"D3",X"13",X"09",X"F3",X"64",X"E3",X"DE",X"C3",X"7C",X"07",X"D6",X"01",X"1A",X"DC",
		X"64",X"C3",X"F9",X"25",X"3A",X"EC",X"64",X"FE",X"00",X"08",X"0D",X"09",X"F4",X"64",X"E3",X"4E",
		X"08",X"E2",X"E5",X"29",X"17",X"11",X"D8",X"40",X"09",X"65",X"08",X"3E",X"01",X"06",X"14",X"E5",
		X"BA",X"17",X"3E",X"03",X"E5",X"1C",X"17",X"C3",X"9C",X"25",X"E5",X"FA",X"0B",X"C3",X"A9",X"25",
		X"E5",X"DA",X"0B",X"C3",X"A9",X"25",X"2A",X"D7",X"64",X"EB",X"F5",X"09",X"00",X"00",X"F5",X"31",
		X"F5",X"7E",X"01",X"F5",X"86",X"02",X"47",X"CE",X"27",X"F5",X"5F",X"02",X"E3",X"38",X"E3",X"38",
		X"E3",X"38",X"E3",X"38",X"F5",X"7E",X"00",X"09",X"1C",X"27",X"E3",X"0F",X"E5",X"95",X"17",X"76",
		X"0B",X"56",X"EB",X"E9",X"40",X"27",X"40",X"27",X"41",X"27",X"61",X"27",X"51",X"27",X"71",X"27",
		X"E1",X"F5",X"7E",X"04",X"90",X"F5",X"5F",X"04",X"E1",X"F5",X"7E",X"04",X"80",X"F5",X"5F",X"04",
		X"E1",X"F5",X"7E",X"03",X"80",X"F5",X"5F",X"03",X"E1",X"F5",X"7E",X"03",X"90",X"F5",X"5F",X"03",
		X"E1",X"2A",X"8C",X"64",X"EB",X"F5",X"09",X"00",X"00",X"F5",X"31",X"EB",X"01",X"00",X"64",X"1F",
		X"3F",X"ED",X"42",X"CD",X"F5",X"7E",X"00",X"09",X"84",X"27",X"E3",X"0F",X"E5",X"95",X"17",X"76",
		X"0B",X"56",X"EB",X"E9",X"54",X"10",X"90",X"27",X"D3",X"27",X"4B",X"10",X"6D",X"10",X"80",X"10",
		X"F5",X"7E",X"03",X"1A",X"8A",X"64",X"F5",X"7E",X"04",X"1A",X"8B",X"64",X"E5",X"EA",X"10",X"F5",
		X"7E",X"06",X"12",X"3A",X"50",X"64",X"FE",X"00",X"08",X"17",X"3A",X"51",X"64",X"FE",X"00",X"08",
		X"17",X"C1",X"09",X"52",X"64",X"21",X"CD",X"D1",X"13",X"01",X"05",X"00",X"1E",X"FF",X"ED",X"98",
		X"E1",X"F5",X"7E",X"06",X"13",X"12",X"30",X"E9",X"F5",X"7E",X"06",X"09",X"08",X"00",X"31",X"EB",
		X"12",X"30",X"F6",X"E5",X"12",X"11",X"F5",X"7E",X"03",X"90",X"1A",X"8A",X"64",X"F5",X"7E",X"04",
		X"1A",X"8B",X"64",X"E5",X"EA",X"10",X"3A",X"50",X"64",X"FE",X"00",X"28",X"1A",X"3A",X"50",X"64",
		X"E3",X"0F",X"F5",X"46",X"05",X"80",X"3D",X"C1",X"FD",X"09",X"52",X"64",X"FD",X"21",X"FD",X"5B");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
